library verilog;
use verilog.vl_types.all;
entity pipelineCycle_vlg_vec_tst is
end pipelineCycle_vlg_vec_tst;
