library verilog;
use verilog.vl_types.all;
entity singleCycle_vlg_vec_tst is
end singleCycle_vlg_vec_tst;
